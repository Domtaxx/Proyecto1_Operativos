// platform.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module platform (
		input  wire        clk_clk,                                  //                               clk.clk
		output wire [12:0] memory_mem_a,                             //                            memory.mem_a
		output wire [2:0]  memory_mem_ba,                            //                                  .mem_ba
		output wire        memory_mem_ck,                            //                                  .mem_ck
		output wire        memory_mem_ck_n,                          //                                  .mem_ck_n
		output wire        memory_mem_cke,                           //                                  .mem_cke
		output wire        memory_mem_cs_n,                          //                                  .mem_cs_n
		output wire        memory_mem_ras_n,                         //                                  .mem_ras_n
		output wire        memory_mem_cas_n,                         //                                  .mem_cas_n
		output wire        memory_mem_we_n,                          //                                  .mem_we_n
		output wire        memory_mem_reset_n,                       //                                  .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,                            //                                  .mem_dq
		inout  wire        memory_mem_dqs,                           //                                  .mem_dqs
		inout  wire        memory_mem_dqs_n,                         //                                  .mem_dqs_n
		output wire        memory_mem_odt,                           //                                  .mem_odt
		output wire        memory_mem_dm,                            //                                  .mem_dm
		input  wire        memory_oct_rzqin,                         //                                  .oct_rzqin
		input  wire        pio_0_external_connection_export,         //         pio_0_external_connection.export
		output wire [6:0]  pio_display_0_external_connection_export, // pio_display_0_external_connection.export
		input  wire [3:0]  pio_password_external_connection_export,  //  pio_password_external_connection.export
		input  wire        rst_reset,                                //                               rst.reset
		output wire        sdram_clk_clk,                            //                         sdram_clk.clk
		output wire [11:0] sdram_wire_addr,                          //                        sdram_wire.addr
		output wire        sdram_wire_ba,                            //                                  .ba
		output wire        sdram_wire_cas_n,                         //                                  .cas_n
		output wire        sdram_wire_cke,                           //                                  .cke
		output wire [3:0]  sdram_wire_cs_n,                          //                                  .cs_n
		inout  wire [63:0] sdram_wire_dq,                            //                                  .dq
		output wire [7:0]  sdram_wire_dqm,                           //                                  .dqm
		output wire        sdram_wire_ras_n,                         //                                  .ras_n
		output wire        sdram_wire_we_n                           //                                  .we_n
	);

	wire         clk_sys_clk_clk;                               // clk:sys_clk_clk -> [HPS:h2f_axi_clk, SDRAM:clk, irq_mapper:clk, mm_interconnect_0:clk_sys_clk_clk, mm_interconnect_1:clk_sys_clk_clk, nios2:clk, pio_0:clk, pio_display_0:clk, pio_password:clk, rom:clk, rst_controller:clk, rst_controller_001:clk]
	wire  [31:0] nios2_data_master_readdata;                    // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_waitrequest;                 // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire  [25:0] nios2_data_master_address;                     // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                  // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire         nios2_data_master_read;                        // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire         nios2_data_master_write;                       // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                   // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire   [1:0] hps_h2f_axi_master_awburst;                    // HPS:h2f_AWBURST -> mm_interconnect_0:HPS_h2f_axi_master_awburst
	wire   [3:0] hps_h2f_axi_master_arlen;                      // HPS:h2f_ARLEN -> mm_interconnect_0:HPS_h2f_axi_master_arlen
	wire   [7:0] hps_h2f_axi_master_wstrb;                      // HPS:h2f_WSTRB -> mm_interconnect_0:HPS_h2f_axi_master_wstrb
	wire         hps_h2f_axi_master_wready;                     // mm_interconnect_0:HPS_h2f_axi_master_wready -> HPS:h2f_WREADY
	wire  [11:0] hps_h2f_axi_master_rid;                        // mm_interconnect_0:HPS_h2f_axi_master_rid -> HPS:h2f_RID
	wire         hps_h2f_axi_master_rready;                     // HPS:h2f_RREADY -> mm_interconnect_0:HPS_h2f_axi_master_rready
	wire   [3:0] hps_h2f_axi_master_awlen;                      // HPS:h2f_AWLEN -> mm_interconnect_0:HPS_h2f_axi_master_awlen
	wire  [11:0] hps_h2f_axi_master_wid;                        // HPS:h2f_WID -> mm_interconnect_0:HPS_h2f_axi_master_wid
	wire   [3:0] hps_h2f_axi_master_arcache;                    // HPS:h2f_ARCACHE -> mm_interconnect_0:HPS_h2f_axi_master_arcache
	wire         hps_h2f_axi_master_wvalid;                     // HPS:h2f_WVALID -> mm_interconnect_0:HPS_h2f_axi_master_wvalid
	wire  [29:0] hps_h2f_axi_master_araddr;                     // HPS:h2f_ARADDR -> mm_interconnect_0:HPS_h2f_axi_master_araddr
	wire   [2:0] hps_h2f_axi_master_arprot;                     // HPS:h2f_ARPROT -> mm_interconnect_0:HPS_h2f_axi_master_arprot
	wire   [2:0] hps_h2f_axi_master_awprot;                     // HPS:h2f_AWPROT -> mm_interconnect_0:HPS_h2f_axi_master_awprot
	wire  [63:0] hps_h2f_axi_master_wdata;                      // HPS:h2f_WDATA -> mm_interconnect_0:HPS_h2f_axi_master_wdata
	wire         hps_h2f_axi_master_arvalid;                    // HPS:h2f_ARVALID -> mm_interconnect_0:HPS_h2f_axi_master_arvalid
	wire   [3:0] hps_h2f_axi_master_awcache;                    // HPS:h2f_AWCACHE -> mm_interconnect_0:HPS_h2f_axi_master_awcache
	wire  [11:0] hps_h2f_axi_master_arid;                       // HPS:h2f_ARID -> mm_interconnect_0:HPS_h2f_axi_master_arid
	wire   [1:0] hps_h2f_axi_master_arlock;                     // HPS:h2f_ARLOCK -> mm_interconnect_0:HPS_h2f_axi_master_arlock
	wire   [1:0] hps_h2f_axi_master_awlock;                     // HPS:h2f_AWLOCK -> mm_interconnect_0:HPS_h2f_axi_master_awlock
	wire  [29:0] hps_h2f_axi_master_awaddr;                     // HPS:h2f_AWADDR -> mm_interconnect_0:HPS_h2f_axi_master_awaddr
	wire   [1:0] hps_h2f_axi_master_bresp;                      // mm_interconnect_0:HPS_h2f_axi_master_bresp -> HPS:h2f_BRESP
	wire         hps_h2f_axi_master_arready;                    // mm_interconnect_0:HPS_h2f_axi_master_arready -> HPS:h2f_ARREADY
	wire  [63:0] hps_h2f_axi_master_rdata;                      // mm_interconnect_0:HPS_h2f_axi_master_rdata -> HPS:h2f_RDATA
	wire         hps_h2f_axi_master_awready;                    // mm_interconnect_0:HPS_h2f_axi_master_awready -> HPS:h2f_AWREADY
	wire   [1:0] hps_h2f_axi_master_arburst;                    // HPS:h2f_ARBURST -> mm_interconnect_0:HPS_h2f_axi_master_arburst
	wire   [2:0] hps_h2f_axi_master_arsize;                     // HPS:h2f_ARSIZE -> mm_interconnect_0:HPS_h2f_axi_master_arsize
	wire         hps_h2f_axi_master_bready;                     // HPS:h2f_BREADY -> mm_interconnect_0:HPS_h2f_axi_master_bready
	wire         hps_h2f_axi_master_rlast;                      // mm_interconnect_0:HPS_h2f_axi_master_rlast -> HPS:h2f_RLAST
	wire         hps_h2f_axi_master_wlast;                      // HPS:h2f_WLAST -> mm_interconnect_0:HPS_h2f_axi_master_wlast
	wire   [1:0] hps_h2f_axi_master_rresp;                      // mm_interconnect_0:HPS_h2f_axi_master_rresp -> HPS:h2f_RRESP
	wire  [11:0] hps_h2f_axi_master_awid;                       // HPS:h2f_AWID -> mm_interconnect_0:HPS_h2f_axi_master_awid
	wire  [11:0] hps_h2f_axi_master_bid;                        // mm_interconnect_0:HPS_h2f_axi_master_bid -> HPS:h2f_BID
	wire         hps_h2f_axi_master_bvalid;                     // mm_interconnect_0:HPS_h2f_axi_master_bvalid -> HPS:h2f_BVALID
	wire   [2:0] hps_h2f_axi_master_awsize;                     // HPS:h2f_AWSIZE -> mm_interconnect_0:HPS_h2f_axi_master_awsize
	wire         hps_h2f_axi_master_awvalid;                    // HPS:h2f_AWVALID -> mm_interconnect_0:HPS_h2f_axi_master_awvalid
	wire         hps_h2f_axi_master_rvalid;                     // mm_interconnect_0:HPS_h2f_axi_master_rvalid -> HPS:h2f_RVALID
	wire         mm_interconnect_0_sdram_s1_chipselect;         // mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	wire  [63:0] mm_interconnect_0_sdram_s1_readdata;           // SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;        // SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	wire  [22:0] mm_interconnect_0_sdram_s1_address;            // mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	wire         mm_interconnect_0_sdram_s1_read;               // mm_interconnect_0:SDRAM_s1_read -> SDRAM:az_rd_n
	wire   [7:0] mm_interconnect_0_sdram_s1_byteenable;         // mm_interconnect_0:SDRAM_s1_byteenable -> SDRAM:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;      // SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;              // mm_interconnect_0:SDRAM_s1_write -> SDRAM:az_wr_n
	wire  [63:0] mm_interconnect_0_sdram_s1_writedata;          // mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	wire         mm_interconnect_0_pio_display_0_s1_chipselect; // mm_interconnect_0:pio_display_0_s1_chipselect -> pio_display_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_display_0_s1_readdata;   // pio_display_0:readdata -> mm_interconnect_0:pio_display_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_display_0_s1_address;    // mm_interconnect_0:pio_display_0_s1_address -> pio_display_0:address
	wire         mm_interconnect_0_pio_display_0_s1_write;      // mm_interconnect_0:pio_display_0_s1_write -> pio_display_0:write_n
	wire  [31:0] mm_interconnect_0_pio_display_0_s1_writedata;  // mm_interconnect_0:pio_display_0_s1_writedata -> pio_display_0:writedata
	wire         mm_interconnect_0_pio_password_s1_chipselect;  // mm_interconnect_0:pio_password_s1_chipselect -> pio_password:chipselect
	wire  [31:0] mm_interconnect_0_pio_password_s1_readdata;    // pio_password:readdata -> mm_interconnect_0:pio_password_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_password_s1_address;     // mm_interconnect_0:pio_password_s1_address -> pio_password:address
	wire         mm_interconnect_0_pio_password_s1_write;       // mm_interconnect_0:pio_password_s1_write -> pio_password:write_n
	wire  [31:0] mm_interconnect_0_pio_password_s1_writedata;   // mm_interconnect_0:pio_password_s1_writedata -> pio_password:writedata
	wire         mm_interconnect_0_pio_0_s1_chipselect;         // mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;           // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_0_s1_address;            // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire         mm_interconnect_0_pio_0_s1_write;              // mm_interconnect_0:pio_0_s1_write -> pio_0:write_n
	wire  [31:0] mm_interconnect_0_pio_0_s1_writedata;          // mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	wire  [31:0] nios2_instruction_master_readdata;             // mm_interconnect_1:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_waitrequest;          // mm_interconnect_1:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [26:0] nios2_instruction_master_address;              // nios2:i_address -> mm_interconnect_1:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                 // nios2:i_read -> mm_interconnect_1:nios2_instruction_master_read
	wire         mm_interconnect_1_rom_s1_chipselect;           // mm_interconnect_1:rom_s1_chipselect -> rom:chipselect
	wire  [31:0] mm_interconnect_1_rom_s1_readdata;             // rom:readdata -> mm_interconnect_1:rom_s1_readdata
	wire         mm_interconnect_1_rom_s1_debugaccess;          // mm_interconnect_1:rom_s1_debugaccess -> rom:debugaccess
	wire  [11:0] mm_interconnect_1_rom_s1_address;              // mm_interconnect_1:rom_s1_address -> rom:address
	wire   [3:0] mm_interconnect_1_rom_s1_byteenable;           // mm_interconnect_1:rom_s1_byteenable -> rom:byteenable
	wire         mm_interconnect_1_rom_s1_write;                // mm_interconnect_1:rom_s1_write -> rom:write
	wire  [31:0] mm_interconnect_1_rom_s1_writedata;            // mm_interconnect_1:rom_s1_writedata -> rom:writedata
	wire         mm_interconnect_1_rom_s1_clken;                // mm_interconnect_1:rom_s1_clken -> rom:clken
	wire         irq_mapper_receiver0_irq;                      // pio_password:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                      // pio_0:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_irq_irq;                                 // irq_mapper:sender_irq -> nios2:irq
	wire         rst_controller_reset_out_reset;                // rst_controller:reset_out -> [SDRAM:reset_n, irq_mapper:reset, mm_interconnect_0:nios2_reset_reset_bridge_in_reset_reset, mm_interconnect_1:nios2_reset_reset_bridge_in_reset_reset, nios2:reset_n, pio_0:reset_n, pio_display_0:reset_n, pio_password:reset_n, rom:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;            // rst_controller:reset_req -> [rom:reset_req, rst_translator:reset_req_in]
	wire         clk_reset_source_reset;                        // clk:reset_source_reset -> rst_controller:reset_in0
	wire         rst_controller_001_reset_out_reset;            // rst_controller_001:reset_out -> mm_interconnect_0:HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	wire         hps_h2f_reset_reset;                           // HPS:h2f_rst_n -> rst_controller_001:reset_in0

	platform_HPS #(
		.F2S_Width (0),
		.S2F_Width (2)
	) hps (
		.mem_a       (memory_mem_a),               //         memory.mem_a
		.mem_ba      (memory_mem_ba),              //               .mem_ba
		.mem_ck      (memory_mem_ck),              //               .mem_ck
		.mem_ck_n    (memory_mem_ck_n),            //               .mem_ck_n
		.mem_cke     (memory_mem_cke),             //               .mem_cke
		.mem_cs_n    (memory_mem_cs_n),            //               .mem_cs_n
		.mem_ras_n   (memory_mem_ras_n),           //               .mem_ras_n
		.mem_cas_n   (memory_mem_cas_n),           //               .mem_cas_n
		.mem_we_n    (memory_mem_we_n),            //               .mem_we_n
		.mem_reset_n (memory_mem_reset_n),         //               .mem_reset_n
		.mem_dq      (memory_mem_dq),              //               .mem_dq
		.mem_dqs     (memory_mem_dqs),             //               .mem_dqs
		.mem_dqs_n   (memory_mem_dqs_n),           //               .mem_dqs_n
		.mem_odt     (memory_mem_odt),             //               .mem_odt
		.mem_dm      (memory_mem_dm),              //               .mem_dm
		.oct_rzqin   (memory_oct_rzqin),           //               .oct_rzqin
		.h2f_rst_n   (hps_h2f_reset_reset),        //      h2f_reset.reset_n
		.h2f_axi_clk (clk_sys_clk_clk),            //  h2f_axi_clock.clk
		.h2f_AWID    (hps_h2f_axi_master_awid),    // h2f_axi_master.awid
		.h2f_AWADDR  (hps_h2f_axi_master_awaddr),  //               .awaddr
		.h2f_AWLEN   (hps_h2f_axi_master_awlen),   //               .awlen
		.h2f_AWSIZE  (hps_h2f_axi_master_awsize),  //               .awsize
		.h2f_AWBURST (hps_h2f_axi_master_awburst), //               .awburst
		.h2f_AWLOCK  (hps_h2f_axi_master_awlock),  //               .awlock
		.h2f_AWCACHE (hps_h2f_axi_master_awcache), //               .awcache
		.h2f_AWPROT  (hps_h2f_axi_master_awprot),  //               .awprot
		.h2f_AWVALID (hps_h2f_axi_master_awvalid), //               .awvalid
		.h2f_AWREADY (hps_h2f_axi_master_awready), //               .awready
		.h2f_WID     (hps_h2f_axi_master_wid),     //               .wid
		.h2f_WDATA   (hps_h2f_axi_master_wdata),   //               .wdata
		.h2f_WSTRB   (hps_h2f_axi_master_wstrb),   //               .wstrb
		.h2f_WLAST   (hps_h2f_axi_master_wlast),   //               .wlast
		.h2f_WVALID  (hps_h2f_axi_master_wvalid),  //               .wvalid
		.h2f_WREADY  (hps_h2f_axi_master_wready),  //               .wready
		.h2f_BID     (hps_h2f_axi_master_bid),     //               .bid
		.h2f_BRESP   (hps_h2f_axi_master_bresp),   //               .bresp
		.h2f_BVALID  (hps_h2f_axi_master_bvalid),  //               .bvalid
		.h2f_BREADY  (hps_h2f_axi_master_bready),  //               .bready
		.h2f_ARID    (hps_h2f_axi_master_arid),    //               .arid
		.h2f_ARADDR  (hps_h2f_axi_master_araddr),  //               .araddr
		.h2f_ARLEN   (hps_h2f_axi_master_arlen),   //               .arlen
		.h2f_ARSIZE  (hps_h2f_axi_master_arsize),  //               .arsize
		.h2f_ARBURST (hps_h2f_axi_master_arburst), //               .arburst
		.h2f_ARLOCK  (hps_h2f_axi_master_arlock),  //               .arlock
		.h2f_ARCACHE (hps_h2f_axi_master_arcache), //               .arcache
		.h2f_ARPROT  (hps_h2f_axi_master_arprot),  //               .arprot
		.h2f_ARVALID (hps_h2f_axi_master_arvalid), //               .arvalid
		.h2f_ARREADY (hps_h2f_axi_master_arready), //               .arready
		.h2f_RID     (hps_h2f_axi_master_rid),     //               .rid
		.h2f_RDATA   (hps_h2f_axi_master_rdata),   //               .rdata
		.h2f_RRESP   (hps_h2f_axi_master_rresp),   //               .rresp
		.h2f_RLAST   (hps_h2f_axi_master_rlast),   //               .rlast
		.h2f_RVALID  (hps_h2f_axi_master_rvalid),  //               .rvalid
		.h2f_RREADY  (hps_h2f_axi_master_rready)   //               .rready
	);

	platform_SDRAM sdram (
		.clk            (clk_sys_clk_clk),                          //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	platform_clk clk (
		.ref_clk_clk        (clk_clk),                //      ref_clk.clk
		.ref_reset_reset    (rst_reset),              //    ref_reset.reset
		.sys_clk_clk        (clk_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),          //    sdram_clk.clk
		.reset_source_reset (clk_reset_source_reset)  // reset_source.reset
	);

	platform_nios2 nios2 (
		.clk           (clk_sys_clk_clk),                      //                       clk.clk
		.reset_n       (~rst_controller_reset_out_reset),      //                     reset.reset_n
		.d_address     (nios2_data_master_address),            //               data_master.address
		.d_byteenable  (nios2_data_master_byteenable),         //                          .byteenable
		.d_read        (nios2_data_master_read),               //                          .read
		.d_readdata    (nios2_data_master_readdata),           //                          .readdata
		.d_waitrequest (nios2_data_master_waitrequest),        //                          .waitrequest
		.d_write       (nios2_data_master_write),              //                          .write
		.d_writedata   (nios2_data_master_writedata),          //                          .writedata
		.i_address     (nios2_instruction_master_address),     //        instruction_master.address
		.i_read        (nios2_instruction_master_read),        //                          .read
		.i_readdata    (nios2_instruction_master_readdata),    //                          .readdata
		.i_waitrequest (nios2_instruction_master_waitrequest), //                          .waitrequest
		.irq           (nios2_irq_irq),                        //                       irq.irq
		.dummy_ci_port ()                                      // custom_instruction_master.readra
	);

	platform_pio_0 pio_0 (
		.clk        (clk_sys_clk_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_0_s1_readdata),   //                    .readdata
		.in_port    (pio_0_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver1_irq)               //                 irq.irq
	);

	platform_pio_display_0 pio_display_0 (
		.clk        (clk_sys_clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_pio_display_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_display_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_display_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_display_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_display_0_s1_readdata),   //                    .readdata
		.out_port   (pio_display_0_external_connection_export)       // external_connection.export
	);

	platform_pio_password pio_password (
		.clk        (clk_sys_clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_pio_password_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_password_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_password_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_password_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_password_s1_readdata),   //                    .readdata
		.in_port    (pio_password_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver0_irq)                      //                 irq.irq
	);

	platform_rom rom (
		.clk         (clk_sys_clk_clk),                      //   clk1.clk
		.address     (mm_interconnect_1_rom_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_1_rom_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_1_rom_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_1_rom_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_1_rom_s1_write),       //       .write
		.readdata    (mm_interconnect_1_rom_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_1_rom_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_1_rom_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze      (1'b0)                                  // (terminated)
	);

	platform_mm_interconnect_0 mm_interconnect_0 (
		.HPS_h2f_axi_master_awid                                        (hps_h2f_axi_master_awid),                       //                                       HPS_h2f_axi_master.awid
		.HPS_h2f_axi_master_awaddr                                      (hps_h2f_axi_master_awaddr),                     //                                                         .awaddr
		.HPS_h2f_axi_master_awlen                                       (hps_h2f_axi_master_awlen),                      //                                                         .awlen
		.HPS_h2f_axi_master_awsize                                      (hps_h2f_axi_master_awsize),                     //                                                         .awsize
		.HPS_h2f_axi_master_awburst                                     (hps_h2f_axi_master_awburst),                    //                                                         .awburst
		.HPS_h2f_axi_master_awlock                                      (hps_h2f_axi_master_awlock),                     //                                                         .awlock
		.HPS_h2f_axi_master_awcache                                     (hps_h2f_axi_master_awcache),                    //                                                         .awcache
		.HPS_h2f_axi_master_awprot                                      (hps_h2f_axi_master_awprot),                     //                                                         .awprot
		.HPS_h2f_axi_master_awvalid                                     (hps_h2f_axi_master_awvalid),                    //                                                         .awvalid
		.HPS_h2f_axi_master_awready                                     (hps_h2f_axi_master_awready),                    //                                                         .awready
		.HPS_h2f_axi_master_wid                                         (hps_h2f_axi_master_wid),                        //                                                         .wid
		.HPS_h2f_axi_master_wdata                                       (hps_h2f_axi_master_wdata),                      //                                                         .wdata
		.HPS_h2f_axi_master_wstrb                                       (hps_h2f_axi_master_wstrb),                      //                                                         .wstrb
		.HPS_h2f_axi_master_wlast                                       (hps_h2f_axi_master_wlast),                      //                                                         .wlast
		.HPS_h2f_axi_master_wvalid                                      (hps_h2f_axi_master_wvalid),                     //                                                         .wvalid
		.HPS_h2f_axi_master_wready                                      (hps_h2f_axi_master_wready),                     //                                                         .wready
		.HPS_h2f_axi_master_bid                                         (hps_h2f_axi_master_bid),                        //                                                         .bid
		.HPS_h2f_axi_master_bresp                                       (hps_h2f_axi_master_bresp),                      //                                                         .bresp
		.HPS_h2f_axi_master_bvalid                                      (hps_h2f_axi_master_bvalid),                     //                                                         .bvalid
		.HPS_h2f_axi_master_bready                                      (hps_h2f_axi_master_bready),                     //                                                         .bready
		.HPS_h2f_axi_master_arid                                        (hps_h2f_axi_master_arid),                       //                                                         .arid
		.HPS_h2f_axi_master_araddr                                      (hps_h2f_axi_master_araddr),                     //                                                         .araddr
		.HPS_h2f_axi_master_arlen                                       (hps_h2f_axi_master_arlen),                      //                                                         .arlen
		.HPS_h2f_axi_master_arsize                                      (hps_h2f_axi_master_arsize),                     //                                                         .arsize
		.HPS_h2f_axi_master_arburst                                     (hps_h2f_axi_master_arburst),                    //                                                         .arburst
		.HPS_h2f_axi_master_arlock                                      (hps_h2f_axi_master_arlock),                     //                                                         .arlock
		.HPS_h2f_axi_master_arcache                                     (hps_h2f_axi_master_arcache),                    //                                                         .arcache
		.HPS_h2f_axi_master_arprot                                      (hps_h2f_axi_master_arprot),                     //                                                         .arprot
		.HPS_h2f_axi_master_arvalid                                     (hps_h2f_axi_master_arvalid),                    //                                                         .arvalid
		.HPS_h2f_axi_master_arready                                     (hps_h2f_axi_master_arready),                    //                                                         .arready
		.HPS_h2f_axi_master_rid                                         (hps_h2f_axi_master_rid),                        //                                                         .rid
		.HPS_h2f_axi_master_rdata                                       (hps_h2f_axi_master_rdata),                      //                                                         .rdata
		.HPS_h2f_axi_master_rresp                                       (hps_h2f_axi_master_rresp),                      //                                                         .rresp
		.HPS_h2f_axi_master_rlast                                       (hps_h2f_axi_master_rlast),                      //                                                         .rlast
		.HPS_h2f_axi_master_rvalid                                      (hps_h2f_axi_master_rvalid),                     //                                                         .rvalid
		.HPS_h2f_axi_master_rready                                      (hps_h2f_axi_master_rready),                     //                                                         .rready
		.clk_sys_clk_clk                                                (clk_sys_clk_clk),                               //                                              clk_sys_clk.clk
		.HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),            // HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.nios2_reset_reset_bridge_in_reset_reset                        (rst_controller_reset_out_reset),                //                        nios2_reset_reset_bridge_in_reset.reset
		.nios2_data_master_address                                      (nios2_data_master_address),                     //                                        nios2_data_master.address
		.nios2_data_master_waitrequest                                  (nios2_data_master_waitrequest),                 //                                                         .waitrequest
		.nios2_data_master_byteenable                                   (nios2_data_master_byteenable),                  //                                                         .byteenable
		.nios2_data_master_read                                         (nios2_data_master_read),                        //                                                         .read
		.nios2_data_master_readdata                                     (nios2_data_master_readdata),                    //                                                         .readdata
		.nios2_data_master_write                                        (nios2_data_master_write),                       //                                                         .write
		.nios2_data_master_writedata                                    (nios2_data_master_writedata),                   //                                                         .writedata
		.pio_0_s1_address                                               (mm_interconnect_0_pio_0_s1_address),            //                                                 pio_0_s1.address
		.pio_0_s1_write                                                 (mm_interconnect_0_pio_0_s1_write),              //                                                         .write
		.pio_0_s1_readdata                                              (mm_interconnect_0_pio_0_s1_readdata),           //                                                         .readdata
		.pio_0_s1_writedata                                             (mm_interconnect_0_pio_0_s1_writedata),          //                                                         .writedata
		.pio_0_s1_chipselect                                            (mm_interconnect_0_pio_0_s1_chipselect),         //                                                         .chipselect
		.pio_display_0_s1_address                                       (mm_interconnect_0_pio_display_0_s1_address),    //                                         pio_display_0_s1.address
		.pio_display_0_s1_write                                         (mm_interconnect_0_pio_display_0_s1_write),      //                                                         .write
		.pio_display_0_s1_readdata                                      (mm_interconnect_0_pio_display_0_s1_readdata),   //                                                         .readdata
		.pio_display_0_s1_writedata                                     (mm_interconnect_0_pio_display_0_s1_writedata),  //                                                         .writedata
		.pio_display_0_s1_chipselect                                    (mm_interconnect_0_pio_display_0_s1_chipselect), //                                                         .chipselect
		.pio_password_s1_address                                        (mm_interconnect_0_pio_password_s1_address),     //                                          pio_password_s1.address
		.pio_password_s1_write                                          (mm_interconnect_0_pio_password_s1_write),       //                                                         .write
		.pio_password_s1_readdata                                       (mm_interconnect_0_pio_password_s1_readdata),    //                                                         .readdata
		.pio_password_s1_writedata                                      (mm_interconnect_0_pio_password_s1_writedata),   //                                                         .writedata
		.pio_password_s1_chipselect                                     (mm_interconnect_0_pio_password_s1_chipselect),  //                                                         .chipselect
		.SDRAM_s1_address                                               (mm_interconnect_0_sdram_s1_address),            //                                                 SDRAM_s1.address
		.SDRAM_s1_write                                                 (mm_interconnect_0_sdram_s1_write),              //                                                         .write
		.SDRAM_s1_read                                                  (mm_interconnect_0_sdram_s1_read),               //                                                         .read
		.SDRAM_s1_readdata                                              (mm_interconnect_0_sdram_s1_readdata),           //                                                         .readdata
		.SDRAM_s1_writedata                                             (mm_interconnect_0_sdram_s1_writedata),          //                                                         .writedata
		.SDRAM_s1_byteenable                                            (mm_interconnect_0_sdram_s1_byteenable),         //                                                         .byteenable
		.SDRAM_s1_readdatavalid                                         (mm_interconnect_0_sdram_s1_readdatavalid),      //                                                         .readdatavalid
		.SDRAM_s1_waitrequest                                           (mm_interconnect_0_sdram_s1_waitrequest),        //                                                         .waitrequest
		.SDRAM_s1_chipselect                                            (mm_interconnect_0_sdram_s1_chipselect)          //                                                         .chipselect
	);

	platform_mm_interconnect_1 mm_interconnect_1 (
		.clk_sys_clk_clk                         (clk_sys_clk_clk),                      //                       clk_sys_clk.clk
		.nios2_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),       // nios2_reset_reset_bridge_in_reset.reset
		.nios2_instruction_master_address        (nios2_instruction_master_address),     //          nios2_instruction_master.address
		.nios2_instruction_master_waitrequest    (nios2_instruction_master_waitrequest), //                                  .waitrequest
		.nios2_instruction_master_read           (nios2_instruction_master_read),        //                                  .read
		.nios2_instruction_master_readdata       (nios2_instruction_master_readdata),    //                                  .readdata
		.rom_s1_address                          (mm_interconnect_1_rom_s1_address),     //                            rom_s1.address
		.rom_s1_write                            (mm_interconnect_1_rom_s1_write),       //                                  .write
		.rom_s1_readdata                         (mm_interconnect_1_rom_s1_readdata),    //                                  .readdata
		.rom_s1_writedata                        (mm_interconnect_1_rom_s1_writedata),   //                                  .writedata
		.rom_s1_byteenable                       (mm_interconnect_1_rom_s1_byteenable),  //                                  .byteenable
		.rom_s1_chipselect                       (mm_interconnect_1_rom_s1_chipselect),  //                                  .chipselect
		.rom_s1_clken                            (mm_interconnect_1_rom_s1_clken),       //                                  .clken
		.rom_s1_debugaccess                      (mm_interconnect_1_rom_s1_debugaccess)  //                                  .debugaccess
	);

	platform_irq_mapper irq_mapper (
		.clk           (clk_sys_clk_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (clk_reset_source_reset),             // reset_in0.reset
		.clk            (clk_sys_clk_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_h2f_reset_reset),               // reset_in0.reset
		.clk            (clk_sys_clk_clk),                    //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
